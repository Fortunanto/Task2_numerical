// 32X32 Iterative Multiplier template
module mult32x32_fast (
    input  logic [31:0] a,        // Input a
    input  logic [31:0] b,        // Input b
    input  logic start,           // Start signal
    output logic [63:0] product,  // Miltiplication product
    output logic valid,           // Operation valid indication

    input  logic clk,             // Clock
    input  logic reset            // Reset
);

// Put your code here
// ------------------


// End of your code

endmodule
